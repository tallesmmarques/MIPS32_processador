library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control is
  port (
    
  );

process(opcode, funct)
begin
	
end process